`ifndef RKV_I2C_QUICK_REG_ACCESS_VIRT_SEQ_SV
`define RKV_I2C_QUICK_REG_ACCESS_VIRT_SEQ_SV
class rkv_i2c_quick_reg_access_virt_seq extends rkv_i2c_base_virtual_sequence;
  
  uvm_status_e status;
	bit [31:0] data;
	
  `uvm_object_utils(rkv_i2c_quick_reg_access_virt_seq)

  function new (string name = "rkv_i2c_quick_reg_access_virt_seq");
    super.new(name);
  endfunction

  virtual task body();
    `uvm_info(get_type_name(), "=====================STARTED=====================", UVM_LOW)
    super.body();
	  
	  
	  
	  rgm.IC_CON.SPEED.set('h3);
	  data = rgm.IC_CON.SPEED.get();
	  `uvm_info("MYDATA", $sformatf("RX_TL readed val : %x", data), UVM_LOW)
	  //`uvm_do(apb_cfg_seq);
//    rgm.RX_TL.set(8'b10101000);
//    //#1ms;
//    rgm.RX_TL.mirror(status);
//	  data = rgm.RX_TL.get();
//	  `uvm_info("MYDATA", $sformatf("RX_TL readed val : %x", data), UVM_LOW)
//    // Attach element sequences below
    `uvm_info(get_type_name(), "=====================FINISHED=====================", UVM_LOW)
  endtask

endclass
`endif // RKV_I2C_QUICK_REG_ACCESS_VIRT_SEQ_SV
