`ifndef I2C_MASTER_TIMEOUT_CG_TEST_SV
`define I2C_MASTER_TIMEOUT_CG_TEST_SV

class i2c_master_timeout_cg_test extends rkv_i2c_base_test;
	`uvm_component_utils(i2c_master_timeout_cg_test)
	function new(string name ="i2c_master_timeout_cg_test", uvm_component parent);
		super.new(name, parent);
	endfunction 
	
	function void build_phase(uvm_phase phase);
		super.build_phase(phase);
    super.cfg.master_scoreboard_enable = 0;
    uvm_config_db#(rkv_i2c_config)::set(this,"env","cfg", super.cfg);
	endfunction
	
	task run_phase(uvm_phase phase);
		i2c_master_timeout_cg_virt_seq seq = i2c_master_timeout_cg_virt_seq::type_id::create("seq");
		`uvm_info("SEQ", "sequence starting", UVM_LOW)
		phase.raise_objection(this);
		seq.start(env.sqr);
		phase.drop_objection(this);
		`uvm_info("SEQ", "sequence finished", UVM_LOW)
	endtask
endclass

`endif


