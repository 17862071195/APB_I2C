
/* Source file "
	/home/verifier/Code_VCS/MyIIC/rkv_i2c_tb/sim/out/obj/partitionlib/_vcs_pc_package__h66j1c/_vcs_pc_package_.v
	", line 1 */
(* VCS_LogicalLibrary = "VCS_PARTCOMP_LIB" *)
config pc__vcs_pc_package__config;
	design pc__vcs_pc_package_;
	cell std liblist DEFAULT;
endconfig
`timescale 1ps/1ps
/* Source file "", line 0 */

(* PARTCOMP_DFT_PKG_WRAPPER = 1 *) 
(* VCS_LogicalLibrary = "VCS_PARTCOMP_LIB" *)

`timescale 1ps/1ps
(* orig_name = "pc__vcs_pc_package_" *)
module pc__vcs_pc_package_;

	initial begin : XmrProcess
	  $$compile_pkg(1, "", "std");
	end
endmodule
