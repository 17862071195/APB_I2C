
`ifndef RKV_I2C_USER_ELEMENT_SEQUENCES_SVH
`define RKV_I2C_USER_ELEMENT_SEQUENCES_SVH
	
	`include "apb_user_address_check_seq.sv"
	`include "apb_user_wait_empty_seq.sv"
	`include "apb_noread_packet_seq.sv"
	`include "apb_user_config_seq.sv"
	`include "apb_write_nocheck_packet_seq.sv"

`endif // RKV_I2C_USER_ELEMENT_SEQUENCES_SVH

